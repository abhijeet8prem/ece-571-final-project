module crc_detection(CrcCor,CrcRem);
  //input clock;
  input logic [15:0]CrcRem;
  output reg [31:0] CrcCor;
  int i;
  wire w1[31:0];

  always_comb
    begin
      case (CrcRem)
        16'b0000000000000001	:	CrcCor=32'h1;	
        16'b0000000000000010	:	CrcCor=32'h2;
        16'b0000000000000100	:	CrcCor=32'h4;
        16'b0000000000001000	:	CrcCor=32'h8;	
        16'b0000000000010000	:	CrcCor=32'h10;
        16'b0000000000100000	:	CrcCor=32'h20;
        16'b0000000001000000	:	CrcCor=32'h40;
        16'b0000000010000000	:	CrcCor=32'h80;
        16'b0000000100000000	:	CrcCor=32'h100;
        16'b0000001000000000	:	CrcCor=32'h200;
        16'b0000010000000000	:	CrcCor=32'h400;
        16'b0000100000000000	:	CrcCor=32'h800;
        16'b0001000000000000	:	CrcCor=32'h1000;
        16'b0010000000000000	:	CrcCor=32'h2000;
        16'b0100000000000000	:	CrcCor=32'h4000;
        16'b1000000000000000	:	CrcCor=32'h8000;
        16'b0001000000100000	:	CrcCor=32'h10000;
        16'b0010000001000010	:	CrcCor=32'h20000;
        16'b0100000010000100	:	CrcCor=32'h40000;
        16'b1000000100001000	:	CrcCor=32'h80000;
        16'b0001001000110001	:	CrcCor=32'h100000;
        16'b0010010001100010	:	CrcCor=32'h200000;
        16'b0100100011000100	:	CrcCor=32'h400000;
        16'b1000000100001000	:	CrcCor=32'h800000;
        16'b0011001100110001	:	CrcCor=32'h1000000;
        16'b0110011001100010	:	CrcCor=32'h2000000;
        16'b1100110011000100	:	CrcCor=32'h4000000;
        16'b1000100110101001	:	CrcCor=32'h8000000;
        16'b0000001101110011	:	CrcCor=32'h10000000;
        16'b0000011011100110	:	CrcCor=32'h20000000;
        16'b0000110111001100	:	CrcCor=32'h40000000;
        16'b0001101110011000	:	CrcCor=32'h80000000;
        default: CrcCor = 32'h0;
      endcase
    end
endmodule
