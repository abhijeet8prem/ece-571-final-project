module Correction(CrcRem, tag, CorVec, CorVec4, iserror);
  input [15:0] CrcRem;
  output logic [31:0] CorVec, CorVec4;
  output logic tag, iserror;
  logic [31:0] CorVec1, CorVec2, CorVec3;
  logic [2:0] hit;

  always_comb
    begin
      if(CrcRem == 0)begin
        iserror = 0;
        $display("No errors were found in the transmitted message");
      end else begin
      case (CrcRem)
        16'b0000000000000001	:	CorVec1 = 32'h00000001;	
        16'b0000000000000010	:	CorVec1 = 32'h00000002;
        16'b0000000000000100	:	CorVec1 = 32'h00000004;
        16'b0000000000001000	:	CorVec1 = 32'h00000008;	
        16'b0000000000010000	:	CorVec1 = 32'h00000010;
        16'b0000000000100000	:	CorVec1 = 32'h00000020;
        16'b0000000001000000	:	CorVec1 = 32'h00000040;
        16'b0000000010000000	:	CorVec1 = 32'h00000080;
        16'b0000000100000000	:	CorVec1 = 32'h00000100;
        16'b0000001000000000	:	CorVec1 = 32'h00000200;
        16'b0000010000000000	:	CorVec1 = 32'h00000400;
        16'b0000100000000000	:	CorVec1 = 32'h00000800;
        16'b0001000000000000	:	CorVec1 = 32'h00001000;
        16'b0010000000000000	:	CorVec1 = 32'h00002000;
        16'b0100000000000000	:	CorVec1 = 32'h00004000;
        16'b1000000000000000	:	CorVec1 = 32'h00008000;
        16'b0001000000100000	:	CorVec1 = 32'h00010000;
        16'b0010000001000010	:	CorVec1 = 32'h00020000;
        16'b0100000010000100	:	CorVec1 = 32'h00040000;
        16'b1000000100001000	:	CorVec1 = 32'h00080000;
        16'b0001001000110001	:	CorVec1 = 32'h00100000;
        16'b0010010001100010	:	CorVec1 = 32'h00200000;
        16'b0100100011000100	:	CorVec1 = 32'h00400000;
        16'b1000000100001000	:	CorVec1 = 32'h00800000;
        16'b0011001100110001	:	CorVec1 = 32'h01000000;
        16'b0110011001100010	:	CorVec1 = 32'h02000000;
        16'b1100110011000100	:	CorVec1 = 32'h04000000;
        16'b1000100110101001	:	CorVec1 = 32'h08000000;
        16'b0000001101110011	:	CorVec1 = 32'h10000000;
        16'b0000011011100110	:	CorVec1 = 32'h20000000;
        16'b0000110111001100	:	CorVec1 = 32'h40000000;
        16'b0001101110011000	:	CorVec1 = 32'h80000000;
        default			:	CorVec1 = 32'h00000000;
      endcase
  
      case(CrcRem)
	16'b0000000000000011    :   CorVec2 = 32'h00000003;	
        16'b0000000000000101    :   CorVec2 = 32'h00000005;	
        16'b0000000000000110    :   CorVec2 = 32'h00000006;	
        16'b0000000000001001    :   CorVec2 = 32'h00000009;	
        16'b0000000000001010    :   CorVec2 = 32'h0000000a;	
        16'b0000000000001100    :   CorVec2 = 32'h0000000c;	
        16'b0000000000010001    :   CorVec2 = 32'h00000011;	
        16'b0000000000010010    :   CorVec2 = 32'h00000012;	
        16'b0000000000010100    :   CorVec2 = 32'h00000014;	
        16'b0000000000011000    :   CorVec2 = 32'h00000018;	
        16'b0000000000100010    :   CorVec2 = 32'h00000022;	
        16'b0000000000100100    :   CorVec2 = 32'h00000024;	
        16'b0000000000101000    :   CorVec2 = 32'h00000028;	
        16'b0000000000110000    :   CorVec2 = 32'h00000030;	
        16'b0000000001000001    :   CorVec2 = 32'h00000041;		
        16'b0000000001000100    :   CorVec2 = 32'h00000044;	
        16'b0000000001001000    :   CorVec2 = 32'h00000048;	
        16'b0000000001010000    :   CorVec2 = 32'h00000050;	
        16'b0000000001100000    :   CorVec2 = 32'h00000060;	
        16'b0000000010000001    :   CorVec2 = 32'h00000081;	
        16'b0000000010000010    :   CorVec2 = 32'h00000082;	
        16'b0000000010001000    :   CorVec2 = 32'h00000088;	
        16'b0000000010010000    :   CorVec2 = 32'h00000090;	
        16'b0000000010100000    :   CorVec2 = 32'h000000a0;	
        16'b0000000011000000    :   CorVec2 = 32'h000000c0;	
        16'b0000000100000001    :   CorVec2 = 32'h00000101;	
        16'b0000000100000010    :   CorVec2 = 32'h00000102;	
        16'b0000000100000100    :   CorVec2 = 32'h00000104;	
        16'b0000000100010000    :   CorVec2 = 32'h00000110;	
        16'b0000000100100000    :   CorVec2 = 32'h00000120;	
        16'b0000000101000000    :   CorVec2 = 32'h00000140;	
        16'b0000000101110011    :   CorVec2 = 32'h10000200;	
        16'b0000000110000000    :   CorVec2 = 32'h00000180;	
        16'b0000001000000001    :   CorVec2 = 32'h00000201;	
        16'b0000001000000010    :   CorVec2 = 32'h00000202;	
        16'b0000001000000100    :   CorVec2 = 32'h00000204;	
        16'b0000001000001000    :   CorVec2 = 32'h00000208;		
        16'b0000001000100000    :   CorVec2 = 32'h00000220;	
        16'b0000001000110001    :   CorVec2 = 32'h00101000;	
        16'b0000001001000000    :   CorVec2 = 32'h00000240;	
        16'b0000001001110011    :   CorVec2 = 32'h10000100;	
        16'b0000001010000000    :   CorVec2 = 32'h00000280;	
        16'b0000001011100110    :   CorVec2 = 32'h20000400;	
        16'b0000001100000000    :   CorVec2 = 32'h00000300;	
        16'b0000001100110011    :   CorVec2 = 32'h10000040;	
        16'b0000001101010011    :   CorVec2 = 32'h10000020;	
        16'b0000001101100011    :   CorVec2 = 32'h10000010;	
        16'b0000001101110001    :   CorVec2 = 32'h10000002;	
        16'b0000001101110010    :   CorVec2 = 32'h10000001;	
        16'b0000001101110111    :   CorVec2 = 32'h10000004;	
        16'b0000001101111011    :   CorVec2 = 32'h10000008;	
        16'b0000001111110011    :   CorVec2 = 32'h10000080;	
        16'b0000010000000001    :   CorVec2 = 32'h00000401;	
        16'b0000010000000010    :   CorVec2 = 32'h00000402;	
        16'b0000010000000100    :   CorVec2 = 32'h00000404;	
        16'b0000010000001000    :   CorVec2 = 32'h00000408;	
        16'b0000010000010000    :   CorVec2 = 32'h00000410;	
        16'b0000010001000000    :   CorVec2 = 32'h00000440;	
        16'b0000010001100010    :   CorVec2 = 32'h00202000;	
        16'b0000010010000000    :   CorVec2 = 32'h00000480;	
        16'b0000010011100110    :   CorVec2 = 32'h20000200;	
        16'b0000010100000000    :   CorVec2 = 32'h00000500;	
        16'b0000010110010101    :   CorVec2 = 32'h30000000;	
        16'b0000010111001100    :   CorVec2 = 32'h40000800;	
        16'b0000011000000000    :   CorVec2 = 32'h00000600;	
        16'b0000011001100110    :   CorVec2 = 32'h20000080;	
        16'b0000011010100110    :   CorVec2 = 32'h20000040;	
        16'b0000011011000110    :   CorVec2 = 32'h20000020;	
        16'b0000011011100010    :   CorVec2 = 32'h20000004;	
        16'b0000011011100100    :   CorVec2 = 32'h20000002;	
        16'b0000011011100111    :   CorVec2 = 32'h20000001;	
        16'b0000011011101110    :   CorVec2 = 32'h20000008;	
        16'b0000011011110110    :   CorVec2 = 32'h20000010;	
        16'b0000011101110011    :   CorVec2 = 32'h10000400;	
        16'b0000011111100110    :   CorVec2 = 32'h20000100;	
        16'b0000100000000001    :   CorVec2 = 32'h00000801;	
        16'b0000100000000010    :   CorVec2 = 32'h00000802;	
        16'b0000100000000100    :   CorVec2 = 32'h00000804;	
        16'b0000100000001000    :   CorVec2 = 32'h00000808;	
        16'b0000100000010000    :   CorVec2 = 32'h00000810;	
        16'b0000100000100000    :   CorVec2 = 32'h00000820;	
        16'b0000100010000000    :   CorVec2 = 32'h00000880;	
        16'b0000100010100001    :   CorVec2 = 32'h08080000;	
        16'b0000100011000100    :   CorVec2 = 32'h00404000;	
        16'b0000100100000000    :   CorVec2 = 32'h00000900;	
        16'b0000100111001100    :   CorVec2 = 32'h40000400;	
        16'b0000101000000000    :   CorVec2 = 32'h00000a00;	
        16'b0000101100101010    :   CorVec2 = 32'h60000000;	
        16'b0000101101110011    :   CorVec2 = 32'h10000800;	
        16'b0000101110011000    :   CorVec2 = 32'h80001000;	
        16'b0000101110111001    :   CorVec2 = 32'h80010000;	
        16'b0000110000000000    :   CorVec2 = 32'h00000c00;	
        16'b0000110011001100    :   CorVec2 = 32'h40000100;	
        16'b0000110101001100    :   CorVec2 = 32'h40000080;	
        16'b0000110110001100    :   CorVec2 = 32'h40000040;	
        16'b0000110111000100    :   CorVec2 = 32'h40000008;	
        16'b0000110111001000    :   CorVec2 = 32'h40000004;	
        16'b0000110111001101    :   CorVec2 = 32'h40000001;	
        16'b0000110111001110    :   CorVec2 = 32'h40000002;	
        16'b0000110111011100    :   CorVec2 = 32'h40000010;	
        16'b0000110111101100    :   CorVec2 = 32'h40000020;	
        16'b0000111010111111    :   CorVec2 = 32'h50000000;	
        16'b0000111011100110    :   CorVec2 = 32'h20000800;	
        16'b0000111111001100    :   CorVec2 = 32'h40000200;	
        16'b0001000000000010    :   CorVec2 = 32'h00001002;	
        16'b0001000000000100    :   CorVec2 = 32'h00001004;	
        16'b0001000000001000    :   CorVec2 = 32'h00001008;	
        16'b0001000000010000    :   CorVec2 = 32'h00001010;	
        16'b0001000000100011    :   CorVec2 = 32'h00010002;	
        16'b0001000000100101    :   CorVec2 = 32'h00010004;	
        16'b0001000000101001    :   CorVec2 = 32'h00010008;	
        16'b0001000001000000    :   CorVec2 = 32'h00001040;	
        16'b0001000001100001    :   CorVec2 = 32'h00010040;		
        16'b0001000010100001    :   CorVec2 = 32'h00010080;	
        16'b0001000100000000    :   CorVec2 = 32'h00001100;	
        16'b0001000100100001    :   CorVec2 = 32'h00010100;	
        16'b0001000101000010    :   CorVec2 = 32'h10100000;	
        16'b0001000110001000    :   CorVec2 = 32'h00808000;	
        16'b0001001000000000    :   CorVec2 = 32'h00001200;	
        16'b0001001000010001    :   CorVec2 = 32'h00100020;		
        16'b0001001000110000    :   CorVec2 = 32'h00100001;	
        16'b0001001000110011    :   CorVec2 = 32'h00100002;	
        16'b0001001000110101    :   CorVec2 = 32'h00100004;	
        16'b0001001000111001    :   CorVec2 = 32'h00100008;	
        16'b0001001001110001    :   CorVec2 = 32'h00100040;	
        16'b0001001010110001    :   CorVec2 = 32'h00100080;	
        16'b0001001101010010    :   CorVec2 = 32'h10010000;		
        16'b0001001110011000    :   CorVec2 = 32'h80000800;	
        16'b0001010000000000    :   CorVec2 = 32'h00001400;	
        16'b0001010000100001    :   CorVec2 = 32'h00010400;	
        16'b0001010011010111    :   CorVec2 = 32'h20100000;	
        16'b0001011000110001    :   CorVec2 = 32'h00100400;	
        16'b0001011001010100    :   CorVec2 = 32'hc0000000;	
        16'b0001011011000111    :   CorVec2 = 32'h20010000;	
        16'b0001011011100110    :   CorVec2 = 32'h20001000;	
        16'b0001011101010011    :   CorVec2 = 32'h01200000;	
        16'b0001100000000000    :   CorVec2 = 32'h00001800;	
        16'b0001100011101011    :   CorVec2 = 32'h90000000;	
        16'b0001100110011000    :   CorVec2 = 32'h80000200;	
        16'b0001101000110001    :   CorVec2 = 32'h00100800;	
        16'b0001101010011000    :   CorVec2 = 32'h80000100;	
        16'b0001101100011000    :   CorVec2 = 32'h80000080;	
        16'b0001101110001000    :   CorVec2 = 32'h80000010;	
        16'b0001101110010000    :   CorVec2 = 32'h80000008;	
        16'b0001101110011001    :   CorVec2 = 32'h80000001;	
        16'b0001101110011010    :   CorVec2 = 32'h80000002;	
        16'b0001101110011100    :   CorVec2 = 32'h80000004;	
        16'b0001101110111000    :   CorVec2 = 32'h80000020;	
        16'b0001101111011000    :   CorVec2 = 32'h80000040;	
        16'b0001110101111110    :   CorVec2 = 32'ha0000000;	
        16'b0001110111001100    :   CorVec2 = 32'h40001000;	
        16'b0001110111101101    :   CorVec2 = 32'h40010000;	
        16'b0001111110011000    :   CorVec2 = 32'h80000400;	
        16'b0001111111111101    :   CorVec2 = 32'h40100000;	
        16'b0010000000000001    :   CorVec2 = 32'h00002001;		
        16'b0010000000000100    :   CorVec2 = 32'h00002004;	
        16'b0010000000001000    :   CorVec2 = 32'h00002008;	
        16'b0010000000010000    :   CorVec2 = 32'h00002010;	
        16'b0010000000100000    :   CorVec2 = 32'h00002020;	
        16'b0010000001000011    :   CorVec2 = 32'h00020001;	
        16'b0010000001000110    :   CorVec2 = 32'h00020004;	
        16'b0010000001001010    :   CorVec2 = 32'h00020008;	
        16'b0010000001010010    :   CorVec2 = 32'h00020010;	
        16'b0010000010000000    :   CorVec2 = 32'h00002080;	
        16'b0010000011000010    :   CorVec2 = 32'h00020080;	
        16'b0010000101000010    :   CorVec2 = 32'h00020100;	
        16'b0010001000000000    :   CorVec2 = 32'h00002200;	
        16'b0010001001000010    :   CorVec2 = 32'h00020200;	
        16'b0010001010000100    :   CorVec2 = 32'h20200000;	
        16'b0010001100010000    :   CorVec2 = 32'h01010000;		
        16'b0010001101110011    :   CorVec2 = 32'h10002000;	
        16'b0010010000000000    :   CorVec2 = 32'h00002400;	
        16'b0010010000100010    :   CorVec2 = 32'h00200040;		
        16'b0010010001100000    :   CorVec2 = 32'h00200002;	
        16'b0010010001100011    :   CorVec2 = 32'h00200001;	
        16'b0010010001100110    :   CorVec2 = 32'h00200004;	
        16'b0010010001101010    :   CorVec2 = 32'h00200008;	
        16'b0010010001110010    :   CorVec2 = 32'h00200010;	
        16'b0010010011100010    :   CorVec2 = 32'h00200080;	
        16'b0010010101100010    :   CorVec2 = 32'h00200100;		
        16'b0010011010100100    :   CorVec2 = 32'h20020000;		
        16'b0010011100010001    :   CorVec2 = 32'h10200000;	
        16'b0010100000000000    :   CorVec2 = 32'h00002800;	
        16'b0010100001000010    :   CorVec2 = 32'h00020800;	
        16'b0010100010101001    :   CorVec2 = 32'h81000000;	
        16'b0010100110101110    :   CorVec2 = 32'h40200000;	
        16'b0010110001100010    :   CorVec2 = 32'h00200800;	
        16'b0010110110001110    :   CorVec2 = 32'h40020000;	
        16'b0010110111001100    :   CorVec2 = 32'h40002000;	
        16'b0010111010100110    :   CorVec2 = 32'h02400000;	
        16'b0011000000000000    :   CorVec2 = 32'h00003000;	
        16'b0011000000100001    :   CorVec2 = 32'h00012000;		
        16'b0011000001100011    :   CorVec2 = 32'h00030000;	
        16'b0011000100110001    :   CorVec2 = 32'h01000200;		
        16'b0011001001110011    :   CorVec2 = 32'h00120000;	
        16'b0011001100010001    :   CorVec2 = 32'h01000020;	
        16'b0011001100100001    :   CorVec2 = 32'h01000010;	
        16'b0011001100110000    :   CorVec2 = 32'h01000001;	
        16'b0011001100110011    :   CorVec2 = 32'h01000002;	
        16'b0011001100110101    :   CorVec2 = 32'h01000004;	
        16'b0011001100111001    :   CorVec2 = 32'h01000008;	
        16'b0011001101110001    :   CorVec2 = 32'h01000040;	
        16'b0011001110110001    :   CorVec2 = 32'h01000080;	
        16'b0011010001000011    :   CorVec2 = 32'h00210000;	
        16'b0011010001100010    :   CorVec2 = 32'h00201000;	
        16'b0011010111010111    :   CorVec2 = 32'h21000000;	
        16'b0011011001010011    :   CorVec2 = 32'h00300000;	
        16'b0011011100110001    :   CorVec2 = 32'h01000400;	
        16'b0011101100110001    :   CorVec2 = 32'h01000800;	
        16'b0011101110011000    :   CorVec2 = 32'h80002000;	
        16'b0011101111011010    :   CorVec2 = 32'h80020000;	
        16'b0011111011111101    :   CorVec2 = 32'h41000000;	
        16'b0011111111111010    :   CorVec2 = 32'h80200000;	
        16'b0100000000000001    :   CorVec2 = 32'h00004001;	
        16'b0100000000000010    :   CorVec2 = 32'h00004002;		
        16'b0100000000001000    :   CorVec2 = 32'h00004008;	
        16'b0100000000010000    :   CorVec2 = 32'h00004010;	
        16'b0100000000100000    :   CorVec2 = 32'h00004020;	
        16'b0100000001000000    :   CorVec2 = 32'h00004040;		
        16'b0100000010000101    :   CorVec2 = 32'h00040001;	
        16'b0100000010000110    :   CorVec2 = 32'h00040002;	
        16'b0100000010001100    :   CorVec2 = 32'h00040008;	
        16'b0100000010010100    :   CorVec2 = 32'h00040010;	
        16'b0100000010100100    :   CorVec2 = 32'h00040020;		
        16'b0100000100000000    :   CorVec2 = 32'h00004100;	
        16'b0100000110000100    :   CorVec2 = 32'h00040100;		
        16'b0100001010000100    :   CorVec2 = 32'h00040200;	
        16'b0100001101110011    :   CorVec2 = 32'h10004000;	
        16'b0100001111110111    :   CorVec2 = 32'h10040000;	
        16'b0100010000000000    :   CorVec2 = 32'h00004400;	
        16'b0100010010000100    :   CorVec2 = 32'h00040400;	
        16'b0100010100001000    :   CorVec2 = 32'h40400000;	
        16'b0100010101101101    :   CorVec2 = 32'h0c000000;	
        16'b0100011000100000    :   CorVec2 = 32'h02020000;	
        16'b0100011011100110    :   CorVec2 = 32'h20004000;	
        16'b0100100000000000    :   CorVec2 = 32'h00004800;	
        16'b0100100001000100    :   CorVec2 = 32'h00400080;	
        16'b0100100011000000    :   CorVec2 = 32'h00400004;	
        16'b0100100011000101    :   CorVec2 = 32'h00400001;	
        16'b0100100011000110    :   CorVec2 = 32'h00400002;	
        16'b0100100011001100    :   CorVec2 = 32'h00400008;	
        16'b0100100011010100    :   CorVec2 = 32'h00400010;	
        16'b0100100011100100    :   CorVec2 = 32'h00400020;	
        16'b0100100111000100    :   CorVec2 = 32'h00400100;	
        16'b0100101011000100    :   CorVec2 = 32'h00400200;	
        16'b0100101110110111    :   CorVec2 = 32'h10400000;		
        16'b0100110101001000    :   CorVec2 = 32'h40040000;	
        16'b0100111000100010    :   CorVec2 = 32'h20400000;	
        16'b0101000000000000    :   CorVec2 = 32'h00005000;	
        16'b0101000000100001    :   CorVec2 = 32'h00014000;	
        16'b0101000010000100    :   CorVec2 = 32'h00041000;	
        16'b0101000010100101    :   CorVec2 = 32'h00050000;	
        16'b0101001000110001    :   CorVec2 = 32'h00104000;	
        16'b0101001010110101    :   CorVec2 = 32'h00140000;	
        16'b0101001101011100    :   CorVec2 = 32'h80400000;	
        16'b0101010101010011    :   CorVec2 = 32'h03000000;	
        16'b0101100011000100    :   CorVec2 = 32'h00401000;	
        16'b0101100011100101    :   CorVec2 = 32'h00410000;	
        16'b0101101011110101    :   CorVec2 = 32'h00500000;	
        16'b0101101100011100    :   CorVec2 = 32'h80040000;	
        16'b0101101110011000    :   CorVec2 = 32'h80004000;	
        16'b0101110101001100    :   CorVec2 = 32'h04800000;	
        16'b0110000000000000    :   CorVec2 = 32'h00006000;	
        16'b0110000001000010    :   CorVec2 = 32'h00024000;		
        16'b0110000011000110    :   CorVec2 = 32'h00060000;	
        16'b0110001001100010    :   CorVec2 = 32'h02000400;		
        16'b0110010011100110    :   CorVec2 = 32'h00240000;	
        16'b0110010100010001    :   CorVec2 = 32'h12000000;	
        16'b0110011000100010    :   CorVec2 = 32'h02000040;	
        16'b0110011001000010    :   CorVec2 = 32'h02000020;	
        16'b0110011001100000    :   CorVec2 = 32'h02000002;	
        16'b0110011001100011    :   CorVec2 = 32'h02000001;	
        16'b0110011001100110    :   CorVec2 = 32'h02000004;	
        16'b0110011001101010    :   CorVec2 = 32'h02000008;	
        16'b0110011001110010    :   CorVec2 = 32'h02000010;	
        16'b0110011011100010    :   CorVec2 = 32'h02000080;	
        16'b0110011101100010    :   CorVec2 = 32'h02000100;	
        16'b0110100010000110    :   CorVec2 = 32'h00420000;	
        16'b0110100011000100    :   CorVec2 = 32'h00402000;	
        16'b0110101110101110    :   CorVec2 = 32'h42000000;	
        16'b0110110010100110    :   CorVec2 = 32'h00600000;	
        16'b0110111001100010    :   CorVec2 = 32'h02000800;	
        16'b0111001100110001    :   CorVec2 = 32'h01004000;	
        16'b0111001110110101    :   CorVec2 = 32'h01040000;	
        16'b0111010001010011    :   CorVec2 = 32'h02100000;	
        16'b0111011001000011    :   CorVec2 = 32'h02010000;	
        16'b0111011001100010    :   CorVec2 = 32'h02001000;	
        16'b0111101111110101    :   CorVec2 = 32'h01400000;	
        16'b0111110111111010    :   CorVec2 = 32'h82000000;	
        16'b1000000000000001    :   CorVec2 = 32'h00008001;	
        16'b1000000000000010    :   CorVec2 = 32'h00008002;	
        16'b1000000000000100    :   CorVec2 = 32'h00008004;		
        16'b1000000000010000    :   CorVec2 = 32'h00008010;	
        16'b1000000000100000    :   CorVec2 = 32'h00008020;	
        16'b1000000001000000    :   CorVec2 = 32'h00008040;	
        16'b1000000010000000    :   CorVec2 = 32'h00008080;	
        16'b1000000100001001    :   CorVec2 = 32'h00080001;	
        16'b1000000100001010    :   CorVec2 = 32'h00080002;	
        16'b1000000100001100    :   CorVec2 = 32'h00080004;	
        16'b1000000100011000    :   CorVec2 = 32'h00080010;	
        16'b1000000100101000    :   CorVec2 = 32'h00080020;	
        16'b1000000101001000    :   CorVec2 = 32'h00080040;		
        16'b1000001000000000    :   CorVec2 = 32'h00008200;	
        16'b1000001001111011    :   CorVec2 = 32'h10080000;	
        16'b1000001100001000    :   CorVec2 = 32'h00080200;	
        16'b1000001101110011    :   CorVec2 = 32'h10008000;	
        16'b1000001110111001    :   CorVec2 = 32'h00900000;	 	
        16'b1000010001100101    :   CorVec2 = 32'h48000000;	
        16'b1000010100001000    :   CorVec2 = 32'h00080400;	
        16'b1000011011100110    :   CorVec2 = 32'h20008000;	
        16'b1000011111101110    :   CorVec2 = 32'h20080000;	
        16'b1000100000000000    :   CorVec2 = 32'h00008800;	
        16'b1000100010101001    :   CorVec2 = 32'h08000100;	
        16'b1000100100001000    :   CorVec2 = 32'h00080800;	
        16'b1000100100101001    :   CorVec2 = 32'h08000080;	
        16'b1000100110001001    :   CorVec2 = 32'h08000020;	
        16'b1000100110100001    :   CorVec2 = 32'h08000008;	
        16'b1000100110101000    :   CorVec2 = 32'h08000001;	
        16'b1000100110101011    :   CorVec2 = 32'h08000002;	
        16'b1000100110101101    :   CorVec2 = 32'h08000004;	
        16'b1000100110111001    :   CorVec2 = 32'h08000010;	
        16'b1000100111101001    :   CorVec2 = 32'h08000040;	
        16'b1000101000010000    :   CorVec2 = 32'h80800000;	
        16'b1000101011011010    :   CorVec2 = 32'h18000000;	
        16'b1000101110101001    :   CorVec2 = 32'h08000200;	
        16'b1000110001000000    :   CorVec2 = 32'h04040000;		
        16'b1000110110101001    :   CorVec2 = 32'h08000400;	
        16'b1000110111001100    :   CorVec2 = 32'h40008000;	
        16'b1000111101001111    :   CorVec2 = 32'h28000000;	
        16'b1001000000000000    :   CorVec2 = 32'h00009000;	
        16'b1001000000100001    :   CorVec2 = 32'h00018000;	
        16'b1001000010001000    :   CorVec2 = 32'h00800100;		
        16'b1001000100101001    :   CorVec2 = 32'h00090000;	
        16'b1001000110000000    :   CorVec2 = 32'h00800008;	
        16'b1001000110001001    :   CorVec2 = 32'h00800001;	
        16'b1001000110001010    :   CorVec2 = 32'h00800002;	
        16'b1001000110001100    :   CorVec2 = 32'h00800004;	
        16'b1001000110011000    :   CorVec2 = 32'h00800010;	
        16'b1001000110101000    :   CorVec2 = 32'h00800020;	
        16'b1001000111001000    :   CorVec2 = 32'h00800040;	
        16'b1001001011111011    :   CorVec2 = 32'h10800000;	
        16'b1001001100111001    :   CorVec2 = 32'h00180000;	
        16'b1001001110001000    :   CorVec2 = 32'h00800200;	
        16'b1001010110001000    :   CorVec2 = 32'h00800400;	
        16'b1001011101101110    :   CorVec2 = 32'h20800000;	
        16'b1001100110101001    :   CorVec2 = 32'h08001000;	
        16'b1001101010010000    :   CorVec2 = 32'h80080000;	
        16'b1001110001000100    :   CorVec2 = 32'h40800000;	
        16'b1010000000000000    :   CorVec2 = 32'h0000a000;	
        16'b1010000001000010    :   CorVec2 = 32'h00028000;	
        16'b1010000100001000    :   CorVec2 = 32'h00082000;	
        16'b1010000101001010    :   CorVec2 = 32'h000a0000;	
        16'b1010001010111001    :   CorVec2 = 32'h01800000;	
        16'b1010010001100010    :   CorVec2 = 32'h00208000;	
        16'b1010010101101010    :   CorVec2 = 32'h00280000;	
        16'b1010100110101001    :   CorVec2 = 32'h08002000;	
        16'b1010100111101011    :   CorVec2 = 32'h08020000;	
        16'b1010101010100110    :   CorVec2 = 32'h06000000;	
        16'b1010110111001011    :   CorVec2 = 32'h08200000;	
        16'b1011000110001000    :   CorVec2 = 32'h00802000;	
        16'b1011000111001010    :   CorVec2 = 32'h00820000;	
        16'b1011001000111001    :   CorVec2 = 32'h01080000;	
        16'b1011001100110001    :   CorVec2 = 32'h01008000;	
        16'b1011010111101010    :   CorVec2 = 32'h00a00000;	
        16'b1011101010011000    :   CorVec2 = 32'h09000000;	
        16'b1100000000000000    :   CorVec2 = 32'h0000c000;	
        16'b1100000010000100    :   CorVec2 = 32'h00048000;	
        16'b1100000101101101    :   CorVec2 = 32'h08400000;	
        16'b1100000110001100    :   CorVec2 = 32'h000c0000;	
        16'b1100010011000100    :   CorVec2 = 32'h04000800;		
        16'b1100100100101101    :   CorVec2 = 32'h08040000;	
        16'b1100100110101001    :   CorVec2 = 32'h08004000;	
        16'b1100100111001100    :   CorVec2 = 32'h00480000;	
        16'b1100101000100010    :   CorVec2 = 32'h24000000;	
        16'b1100110001000100    :   CorVec2 = 32'h04000080;	
        16'b1100110010000100    :   CorVec2 = 32'h04000040;	
        16'b1100110011000000    :   CorVec2 = 32'h04000004;	
        16'b1100110011000101    :   CorVec2 = 32'h04000001;	
        16'b1100110011000110    :   CorVec2 = 32'h04000002;	
        16'b1100110011001100    :   CorVec2 = 32'h04000008;	
        16'b1100110011010100    :   CorVec2 = 32'h04000010;	
        16'b1100110011100100    :   CorVec2 = 32'h04000020;	
        16'b1100110111000100    :   CorVec2 = 32'h04000100;	
        16'b1100111011000100    :   CorVec2 = 32'h04000200;	
        16'b1100111110110111    :   CorVec2 = 32'h14000000;	
        16'b1101000100001100    :   CorVec2 = 32'h00840000;	
        16'b1101000110001000    :   CorVec2 = 32'h00804000;	
        16'b1101011101011100    :   CorVec2 = 32'h84000000;	
        16'b1101100101001100    :   CorVec2 = 32'h00c00000;	
        16'b1101110011000100    :   CorVec2 = 32'h04001000;	
        16'b1101110011100101    :   CorVec2 = 32'h04010000;	
        16'b1101111011110101    :   CorVec2 = 32'h04100000;	
        16'b1110011001100010    :   CorVec2 = 32'h02008000;	
        16'b1110011101101010    :   CorVec2 = 32'h02080000;	
        16'b1110100010100110    :   CorVec2 = 32'h04200000;	
        16'b1110110010000110    :   CorVec2 = 32'h04020000;	
        16'b1110110011000100    :   CorVec2 = 32'h04002000;	
        16'b1110111111001011    :   CorVec2 = 32'h0a000000;	
        16'b1111011111101010    :   CorVec2 = 32'h02800000;	
        16'b1111111111110101    :   CorVec2 = 32'h05000000;	
        default                 :       CorVec2 = 32'h00000000;
      endcase
 
      case(CrcRem)
  	16'b0000000000100001    :       begin
                                        CorVec3 = 32'h00000021;
                                        CorVec4 = 32'h00011000;
                                        end
        16'b0000000001000010    :       begin
                                        CorVec3 = 32'h00000042;
                                        CorVec4 = 32'h00022000;
                                        end
        16'b0000000010000100    :       begin
                                        CorVec3 = 32'h00000084;
                                        CorVec4 = 32'h00044000;
                                        end
        16'b0000000100001000    :       begin
                                        CorVec3 = 32'h00000108;
                                        CorVec4 = 32'h00088000;
                                        end
        16'b0000001000010000    :       begin
                                        CorVec3 = 32'h00000210;
                                        CorVec4 = 32'h00110000;
                                        end
        16'b0000010000100000    :       begin
                                        CorVec3 = 32'h00000420;
                                        CorVec4 = 32'h00220000;
                                        end
        16'b0000100001000000    :       begin
                                        CorVec3 = 32'h00000840;
                                        CorVec4 = 32'h00440000;
                                        end
        16'b0000100110101001    :       begin
                                        CorVec3 = 32'h08008000;
                                        CorVec4 = 32'h80100000;
                                        end
        16'b0001000000000001    :       begin
                                        CorVec3 = 32'h00001001;
                                        CorVec4 = 32'h00010020;
                                        end
        16'b0001000000100000    :       begin
                                        CorVec3 = 32'h00001020;
                                        CorVec4 = 32'h00010001;
                                        end
        16'b0001000000110001    :       begin
                                        CorVec3 = 32'h00010010;
                                        CorVec4 = 32'h00100200;
                                        end
        16'b0001000010000000    :       begin
                                        CorVec3 = 32'h00001080;
                                        CorVec4 = 32'h00880000;
                                        end
        16'b0001001000100001    :       begin
                                        CorVec3 = 32'h00010200;
                                        CorVec4 = 32'h00100010;
                                        end
        16'b0001001100110001    :       begin
                                        CorVec3 = 32'h00100100;
                                        CorVec4 = 32'h01002000;
                                        end
        16'b0001001101110011    :       begin
                                        CorVec3 = 32'h01020000;
                                        CorVec4 = 32'h10001000;
                                        end
        16'b0001100000100001    :       begin
                                        CorVec3 = 32'h00010800;
                                        CorVec4 = 32'h08800000;
                                        end
        16'b0010000000000010    :       begin
                                        CorVec3 = 32'h00002002;
                                        CorVec4 = 32'h00020040;
                                        end
        16'b0010000001000000    :       begin
                                        CorVec3 = 32'h00002040;
                                        CorVec4 = 32'h00020002;
                                        end
        16'b0010000001100010    :       begin
                                        CorVec3 = 32'h00020020;
                                        CorVec4 = 32'h00200400;
                                        end
        16'b0010000100000000    :       begin
                                        CorVec3 = 32'h00002100;
                                        CorVec4 = 32'h01100000;
                                        end
        16'b0010001100110001    :       begin
                                        CorVec3 = 32'h01001000;
                                        CorVec4 = 32'h10020000;
                                        end
        16'b0010010001000010    :       begin 
                                        CorVec3 = 32'h00020400;
                                        CorVec4 = 32'h00200020;
                                        end
        16'b0010011001100010    :       begin 
                                        CorVec3 = 32'h00200200;
                                        CorVec4 = 32'h02004000;
                                        end
        16'b0010011011100110    :       begin 
                                        CorVec3 = 32'h02040000;
                                        CorVec4 = 32'h20002000; 
                                        end
        16'b0011000001000010    :       begin 
                                        CorVec3 = 32'h00021000;
                                        CorVec4 = 32'h11000000;
                                        end
        16'b0011001000110001    :       begin 
                                        CorVec3 = 32'h00102000;
                                        CorVec4 = 32'h01000100;
                                        end
        16'b0100000000000100    :       begin 
                                        CorVec3 = 32'h00004004;
                                        CorVec4 = 32'h00040080;
                                        end
        16'b0100000010000000    :       begin
                                        CorVec3 = 32'h00004080;
                                        CorVec4 = 32'h00040004;
                                        end
        16'b0100000011000100    :       begin 
                                        CorVec3 = 32'h00040040;
                                        CorVec4 = 32'h00400800;
                                        end
        16'b0100001000000000    :       begin 
                                        CorVec3 = 32'h00004200;
                                        CorVec4 = 32'h02200000;
                                        end
        16'b0100011001100010    :       begin 
                                        CorVec3 = 32'h02002000;
                                        CorVec4 = 32'h20040000;
                                        end
        16'b0100100010000100    :       begin
                                        CorVec3 = 32'h00040800;
                                        CorVec4 = 32'h00400040;
                                        end
        16'b0100110011000100    :       begin 
                                        CorVec3 = 32'h00400400;
                                        CorVec4 = 32'h04008000;
                                        end
        16'b0100110111001100    :       begin 
                                        CorVec3 = 32'h04080000;
                                        CorVec4 = 32'h40004000;
                                        end
        16'b0110000010000100    :       begin
                                        CorVec3 = 32'h00042000;
                                        CorVec4 = 32'h22000000;
                                        end 
        16'b0110010001100010    :       begin 
                                        CorVec3 = 32'h00204000;
                                        CorVec4 = 32'h02000200;
                                        end
        16'b1000000000001000    :       begin 
                                        CorVec3 = 32'h00008008;
                                        CorVec4 = 32'h00080100;
                                        end
        16'b1000000100000000    :       begin 
                                        CorVec3 = 32'h00008100;
                                        CorVec4 = 32'h00080008;
                                        end
        16'b1000000110001000    :       begin 
                                        CorVec3 = 32'h00080080;
                                        CorVec4 = 32'h00801000;
                                        end
        16'b1000000110101001    :       begin 
                                        CorVec3 = 32'h00810000;
                                        CorVec4 = 32'h08000800;
                                        end
        16'b1000010000000000    :       begin 
                                        CorVec3 = 32'h00008400;
                                        CorVec4 = 32'h04400000;
                                        end
        16'b1000110011000100    :       begin 
                                        CorVec3 = 32'h04004000;
                                        CorVec4 = 32'h40080000;
                                        end
        16'b1001000100001000    :       begin 
                                        CorVec3 = 32'h00081000;
                                        CorVec4 = 32'h00800080;
                                        end
        16'b1001001000110001    :       begin  
                                        CorVec3 = 32'h00108000;
                                        CorVec4 = 32'h88000000;
                                        end
        16'b1001100110001000    :       begin 
                                        CorVec3 = 32'h00800800;
                                        CorVec4 = 32'h08010000;
                                        end
        16'b1001101110011000    :       begin 
                                        CorVec3 = 32'h08100000;
                                        CorVec4 = 32'h80008000;
                                        end
        16'b1100000100001000    :       begin 
                                        CorVec3 = 32'h00084000;
                                        CorVec4 = 32'h44000000;
                                        end
        16'b1100100011000101    :       begin 
                                        CorVec3 = 32'h00408000;
                                        CorVec4 = 32'h04000400;
                                        end
        default                 :	begin 
					CorVec3 = 32'h00000000;
					CorVec4 = 32'h00000000;
					end
      endcase
      end
    end
  
  always_comb
    begin
      if(CorVec1)
        hit = 3'b100;
      else if(CorVec2)
        hit = 3'b010;
      else if(CorVec3)
        hit = 3'b001;
      else
        hit= 3'b000;
    end
  
  always_comb
    begin
      case(hit)
          3'b100 	: CorVec = CorVec1;
          3'b010 	: CorVec = CorVec2;
          3'b001 	: CorVec = CorVec3;
          default 	: CorVec = '0;
      endcase
    end

endmodule

